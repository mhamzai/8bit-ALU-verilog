module testbench();
reg[3:0] a1,b1;
reg[4:0] switch;
reg cary;
wire [4:0] out;
ALU unit(out,a1,b1,switch,cary);
initial begin
a1[0]=0;
a1[1]=1;
a1[2]=1;
a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=0;
switch[1]=0;
switch[2]=0;
switch[3]=0;
switch[4]=0;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=1;
switch[0]=0;
switch[1]=0;
switch[2]=0;
switch[3]=0;
switch[4]=0;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=0;
switch[1]=1;
switch[2]=0;
switch[3]=0;
switch[4]=0;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=1;
switch[1]=0;
switch[2]=0;
switch[3]=0;
switch[4]=0;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=1;
switch[1]=1;
switch[2]=0;
switch[3]=0;
switch[4]=0;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=0;
switch[1]=0;
switch[2]=0;
switch[3]=0;
switch[4]=1;
#100

a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=0;
switch[1]=0;
switch[2]=0;
switch[3]=1;
switch[4]=1;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=0;
switch[0]=0;
switch[1]=0;
switch[2]=1;
switch[3]=0;
switch[4]=1;
#100
a1[0]=1;a1[1]=1;a1[2]=1;a1[3]=0;
b1[0]=1;b1[1]=0;b1[2]=1;b1[3]=0;
cary=1;
switch[0]=0;
switch[1]=0;
switch[2]=1;
switch[3]=1;
switch[4]=1;
end
endmodule
